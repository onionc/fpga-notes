
`timescale 1 ns / 100 ps
module pic_ram (address, q);

    input wire [8:0] address;
    output reg [800<<2:0] q;
	 
	always @ (*)
		case(address)
			9'd0  : q = 3200'hB93C73448D6C6A7C697CA87C8774667C48842A844984688448844884297C297C497C48844884287C287C087C087C087C087C277C277C267C247CE583C78B0974296C4674257C0784C7734A7C2964EC2B161D950CB424552C333CC9534784C67BEB73B05B53533563D67A948AB28A137B3473F482D482F47A33733373137B3383F26A535BB353934B934BB453B4537453744B744B745374539453945374539453945374535453345B3463546354635463545B545B545B745374537453745374537453545B545B545B545B545B545B545B545B545B545B545B54535453545B555B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B555B555B555B555B555B555B556355635563556355635563556355635563556355635563556355637563745B755B745B745B745B755B565B76639563946395639663935BAC5B8B6C8B6C4A6C8A6C896C686C47648D74B1639663986BD76BD063AA64C8648B5C325C3964D95B;
			9'd1  : q = 3200'hB93C73448D6C6A7C697CA87C8774667C48842A844984688448844884297C297C497C48844884287C287C087C087C087C087C277C277C267C247CE583C78B0974296C4674257C0784C7734A7C2964EC2B161D950CB424552C333CC9534784C67BEB73B05B53533563D67A948AB28A137B3473F482D482F47A33733373137B3383F26A535BB353934B934BB453B4537453744B744B745374539453945374539453945374535453345B3463546354635463545B545B545B745374537453745374537453545B545B545B545B545B545B545B545B545B545B545B54535453545B555B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B555B555B555B555B555B555B556355635563556355635563556355635563556355635563556355637563745B755B745B745B745B755B565B76639563946395639663935BAC5B8B6C8B6C4A6C8A6C896C686C47648D74B1639663986BD76BD063AA64C8648B5C325C3964D95B;
			9'd2  : q = 3200'hB93C73448D6C6A7C697CA87C8774667C48842A844984688448844884297C297C497C48844884287C287C087C087C087C087C277C277C267C247CE583C78B0974296C4674257C0784C7734A7C2964EC2B161D950CB424552C333CC9534784C67BEB73B05B53533563D67A948AB28A137B3473F482D482F47A33733373137B3383F26A535BB353934B934BB453B4537453744B744B745374539453945374539453945374535453345B3463546354635463545B545B545B745374537453745374537453545B545B545B545B545B545B545B545B545B545B545B54535453545B555B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B555B555B555B555B555B555B556355635563556355635563556355635563556355635563556355637563745B755B745B745B745B755B565B76639563946395639663935BAC5B8B6C8B6C4A6C8A6C896C686C47648D74B1639663986BD76BD063AA64C8648B5C325C3964D95B;
			9'd3  : q = 3200'hB93C73448D6C6A7C697CA87C8774667C48842A844984688448844884297C297C497C48844884287C287C087C087C087C087C277C277C267C247CE583C78B0974296C4674257C0784C7734A7C2964EC2B161D950CB424552C333CC9534784C67BEB73B05B53533563D67A948AB28A137B3473F482D482F47A33733373137B3383F26A535BB353934B934BB453B4537453744B744B745374539453945374539453945374535453345B3463546354635463545B545B545B745374537453745374537453545B545B545B545B545B545B545B545B545B545B545B54535453545B555B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B555B555B555B555B555B555B556355635563556355635563556355635563556355635563556355637563745B755B745B745B745B755B565B76639563946395639663935BAC5B8B6C8B6C4A6C8A6C896C686C47648D74B1639663986BD76BD063AA64C8648B5C325C3964D95B;
			9'd4  : q = 3200'hB93C73448D6C6A7C697CA87C8774667C48842A844984688448844884297C297C497C48844884287C287C087C087C087C087C277C277C267C247CE583C78B0974296C4674257C0784C7734A7C2964EC2B161D950CB424552C333CC9534784C67BEB73B05B53533563D67A948AB28A137B3473F482D482F47A33733373137B3383F26A535BB353934B934BB453B4537453744B744B745374539453945374539453945374535453345B3463546354635463545B545B545B745374537453745374537453545B545B545B545B545B545B545B545B545B545B545B54535453545B555B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B555B555B555B555B555B555B556355635563556355635563556355635563556355635563556355637563745B755B745B745B745B755B565B76639563946395639663935BAC5B8B6C8B6C4A6C8A6C896C686C47648D74B1639663986BD76BD063AA64C8648B5C325C3964D95B;
			9'd5  : q = 3200'hB93C73448D6C6A7C697CA87C8774667C48842A844984688448844884297C297C497C48844884287C287C087C087C087C087C277C277C267C247CE583C78B0974296C4674257C0784C7734A7C2964EC2B161D950CB424552C333CC9534784C67BEB73B05B53533563D67A948AB28A137B3473F482D482F47A33733373137B3383F26A535BB353934B934BB453B4537453744B744B745374539453945374539453945374535453345B3463546354635463545B545B545B745374537453745374537453545B545B545B545B545B545B545B545B545B545B545B54535453545B555B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B555B555B555B555B555B555B556355635563556355635563556355635563556355635563556355637563745B755B745B745B745B755B565B76639563946395639663935BAC5B8B6C8B6C4A6C8A6C896C686C47648D74B1639663986BD76BD063AA64C8648B5C325C3964D95B;
			9'd6  : q = 3200'hB93C73448D6C6A7C697CA87C8774667C48842A844984688448844884297C297C497C48844884287C287C087C087C087C087C277C277C267C247CE583C78B0974296C4674257C0784C7734A7C2964EC2B161D950CB424552C333CC9534784C67BEB73B05B53533563D67A948AB28A137B3473F482D482F47A33733373137B3383F26A535BB353934B934BB453B4537453744B744B745374539453945374539453945374535453345B3463546354635463545B545B545B745374537453745374537453545B545B545B545B545B545B545B545B545B545B545B54535453545B555B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B555B555B555B555B555B555B556355635563556355635563556355635563556355635563556355637563745B755B745B745B745B755B565B76639563946395639663935BAC5B8B6C8B6C4A6C8A6C896C686C47648D74B1639663986BD76BD063AA64C8648B5C325C3964D95B;
			9'd7  : q = 3200'hB93C73448D6C6A7C697CA87C8774667C48842A844984688448844884297C297C497C48844884287C287C087C087C087C087C277C277C267C247CE583C78B0974296C4674257C0784C7734A7C2964EC2B161D950CB424552C333CC9534784C67BEB73B05B53533563D67A948AB28A137B3473F482D482F47A33733373137B3383F26A535BB353934B934BB453B4537453744B744B745374539453945374539453945374535453345B3463546354635463545B545B545B745374537453745374537453545B545B545B545B545B545B545B545B545B545B545B54535453545B555B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B555B555B555B555B555B555B556355635563556355635563556355635563556355635563556355637563745B755B745B745B745B755B565B76639563946395639663935BAC5B8B6C8B6C4A6C8A6C896C686C47648D74B1639663986BD76BD063AA64C8648B5C325C3964D95B;
			9'd8  : q = 3200'hB93C73448D6C6A7C697CA87C8774667C48842A844984688448844884297C297C497C48844884287C287C087C087C087C087C277C277C267C247CE583C78B0974296C4674257C0784C7734A7C2964EC2B161D950CB424552C333CC9534784C67BEB73B05B53533563D67A948AB28A137B3473F482D482F47A33733373137B3383F26A535BB353934B934BB453B4537453744B744B745374539453945374539453945374535453345B3463546354635463545B545B545B745374537453745374537453545B545B545B545B545B545B545B545B545B545B545B54535453545B555B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B555B555B555B555B555B555B556355635563556355635563556355635563556355635563556355637563745B755B745B745B745B755B565B76639563946395639663935BAC5B8B6C8B6C4A6C8A6C896C686C47648D74B1639663986BD76BD063AA64C8648B5C325C3964D95B;
			9'd9  : q = 2300'hB93C73448D6C6A7C697CA87C8774667C48842A844984688448844884297C297C497C48844884287C287C087C087C087C087C277C277C267C247CE583C78B0974296C4674257C0784C7734A7C2964EC2B161D950CB424552C333CC9534784C67BEB73B05B53533563D67A948AB28A137B3473F482D482F47A33733373137B3383F26A535BB353934B934BB453B4537453744B744B745374539453945374539453945374535453345B3463546354635463545B545B545B745374537453745374537453545B545B545B545B545B545B545B545B545B545B545B54535453545B555B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B555B555B555B555B555B555B556355635563556355635563556355635563556355635563556355637563745B755B745B745B745B755B565B76639563946395639663935BAC5B8B6C8B6C4A6C8A6C896C686C47648D74B1639663986BD76BD063AA64C8648B5C325C3964D95B;
			//9'd10  : q = 3200'hB93C73448D6C6A7C697CA87C8774667C48842A844984688448844884297C297C497C48844884287C287C087C087C087C087C277C277C267C247CE583C78B0974296C4674257C0784C7734A7C2964EC2B161D950CB424552C333CC9534784C67BEB73B05B53533563D67A948AB28A137B3473F482D482F47A33733373137B3383F26A535BB353934B934BB453B4537453744B744B745374539453945374539453945374535453345B3463546354635463545B545B545B745374537453745374537453545B545B545B545B545B545B545B545B545B545B545B54535453545B555B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B355B555B555B555B555B555B555B556355635563556355635563556355635563556355635563556355637563745B755B745B745B745B755B565B76639563946395639663935BAC5B8B6C8B6C4A6C8A6C896C686C47648D74B1639663986BD76BD063AA64C8648B5C325C3964D95B;
			
			default:q = 0;
			
			
			
		endcase
		
endmodule
